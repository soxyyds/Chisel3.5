module ALU(
  input         clock,
  input         reset,
  input  [31:0] io_src1_in,
  input  [31:0] io_src2_in,
  input  [5:0]  io_instr_id,
  input         io_valid_in,
  input         io_flush_in,
  input  [31:0] io_pc_in,
  input  [31:0] io_imm_in,
  output [31:0] io_result_out,
  output        io_valid_out,
  output        io_branch_out,
  output [31:0] io_jump_addr,
  output        io_is_load,
  output        io_is_store
);
  wire [31:0] _next_pc_T_1 = io_pc_in + 32'h4; // @[ALU.scala 82:23]
  wire [31:0] _result_T_1 = io_src1_in + io_src2_in; // @[ALU.scala 89:38]
  wire [31:0] _result_T_3 = io_src1_in + io_imm_in; // @[ALU.scala 90:38]
  wire [31:0] _result_T_5 = io_src1_in - io_src2_in; // @[ALU.scala 91:38]
  wire [31:0] _result_T_7 = io_pc_in + io_imm_in; // @[ALU.scala 93:36]
  wire [62:0] _GEN_1 = {{31'd0}, io_src1_in}; // @[ALU.scala 94:38]
  wire [62:0] _result_T_9 = _GEN_1 << io_src2_in[4:0]; // @[ALU.scala 94:38]
  wire [62:0] _GEN_3 = {{31'd0}, io_src1_in}; // @[ALU.scala 95:38]
  wire [62:0] _result_T_11 = _GEN_3 << io_imm_in[4:0]; // @[ALU.scala 95:38]
  wire [31:0] _result_T_13 = io_src1_in >> io_src2_in[4:0]; // @[ALU.scala 96:38]
  wire [31:0] _result_T_15 = io_src1_in >> io_imm_in[4:0]; // @[ALU.scala 97:38]
  wire [31:0] _result_T_16 = io_src1_in; // @[ALU.scala 98:39]
  wire [31:0] _result_T_19 = $signed(io_src1_in) >>> io_src2_in[4:0]; // @[ALU.scala 98:67]
  wire [31:0] _result_T_23 = $signed(io_src1_in) >>> io_imm_in[4:0]; // @[ALU.scala 99:66]
  wire [31:0] _result_T_24 = io_src1_in | io_src2_in; // @[ALU.scala 100:38]
  wire [31:0] _result_T_25 = io_src1_in | io_imm_in; // @[ALU.scala 101:38]
  wire [31:0] _result_T_26 = io_src1_in & io_src2_in; // @[ALU.scala 102:38]
  wire [31:0] _result_T_27 = io_src1_in & io_imm_in; // @[ALU.scala 103:38]
  wire [31:0] _result_T_28 = io_src1_in ^ io_src2_in; // @[ALU.scala 104:38]
  wire [31:0] _result_T_29 = io_src1_in ^ io_imm_in; // @[ALU.scala 105:38]
  wire [31:0] _result_T_31 = io_src2_in; // @[ALU.scala 106:59]
  wire  _result_T_32 = $signed(io_src1_in) < $signed(io_src2_in); // @[ALU.scala 106:46]
  wire [31:0] _result_T_34 = io_imm_in; // @[ALU.scala 107:58]
  wire  _result_T_36 = io_src1_in < io_src2_in; // @[ALU.scala 108:39]
  wire [31:0] _next_pc_T_6 = _result_T_3 & 32'hfffffffe; // @[ALU.scala 119:43]
  wire  _GEN_5 = 6'h1c == io_instr_id & io_src1_in >= io_src2_in; // @[ALU.scala 145:20 81:16 87:23]
  wire  _GEN_10 = 6'h1b == io_instr_id ? _result_T_36 : _GEN_5; // @[ALU.scala 141:20 87:23]
  wire  _GEN_15 = 6'h1a == io_instr_id ? $signed(io_src1_in) >= $signed(io_src2_in) : _GEN_10; // @[ALU.scala 137:20 87:23]
  wire  _GEN_20 = 6'h19 == io_instr_id ? _result_T_32 : _GEN_15; // @[ALU.scala 133:20 87:23]
  wire  _GEN_25 = 6'h18 == io_instr_id ? io_src1_in != io_src2_in : _GEN_20; // @[ALU.scala 129:20 87:23]
  wire  _GEN_30 = 6'h17 == io_instr_id ? io_src1_in == io_src2_in : _GEN_25; // @[ALU.scala 125:20 87:23]
  wire  _GEN_37 = 6'h16 == io_instr_id | _GEN_30; // @[ALU.scala 120:20 87:23]
  wire  _GEN_42 = 6'h15 == io_instr_id | _GEN_37; // @[ALU.scala 115:20 87:23]
  wire  _GEN_47 = 6'h14 == io_instr_id ? 1'h0 : _GEN_42; // @[ALU.scala 81:16 87:23]
  wire  _GEN_52 = 6'h13 == io_instr_id ? 1'h0 : _GEN_47; // @[ALU.scala 81:16 87:23]
  wire  _GEN_57 = 6'h12 == io_instr_id ? 1'h0 : _GEN_52; // @[ALU.scala 81:16 87:23]
  wire  _GEN_62 = 6'h11 == io_instr_id ? 1'h0 : _GEN_57; // @[ALU.scala 81:16 87:23]
  wire  _GEN_67 = 6'h10 == io_instr_id ? 1'h0 : _GEN_62; // @[ALU.scala 81:16 87:23]
  wire  _GEN_72 = 6'hf == io_instr_id ? 1'h0 : _GEN_67; // @[ALU.scala 81:16 87:23]
  wire  _GEN_77 = 6'he == io_instr_id ? 1'h0 : _GEN_72; // @[ALU.scala 81:16 87:23]
  wire  _GEN_82 = 6'hd == io_instr_id ? 1'h0 : _GEN_77; // @[ALU.scala 81:16 87:23]
  wire  _GEN_87 = 6'hc == io_instr_id ? 1'h0 : _GEN_82; // @[ALU.scala 81:16 87:23]
  wire  _GEN_92 = 6'hb == io_instr_id ? 1'h0 : _GEN_87; // @[ALU.scala 81:16 87:23]
  wire  _GEN_97 = 6'ha == io_instr_id ? 1'h0 : _GEN_92; // @[ALU.scala 81:16 87:23]
  wire  _GEN_102 = 6'h9 == io_instr_id ? 1'h0 : _GEN_97; // @[ALU.scala 81:16 87:23]
  wire  _GEN_107 = 6'h8 == io_instr_id ? 1'h0 : _GEN_102; // @[ALU.scala 81:16 87:23]
  wire  _GEN_112 = 6'h7 == io_instr_id ? 1'h0 : _GEN_107; // @[ALU.scala 81:16 87:23]
  wire  _GEN_117 = 6'h6 == io_instr_id ? 1'h0 : _GEN_112; // @[ALU.scala 81:16 87:23]
  wire  _GEN_122 = 6'h5 == io_instr_id ? 1'h0 : _GEN_117; // @[ALU.scala 81:16 87:23]
  wire  _GEN_127 = 6'h4 == io_instr_id ? 1'h0 : _GEN_122; // @[ALU.scala 81:16 87:23]
  wire  _GEN_132 = 6'h3 == io_instr_id ? 1'h0 : _GEN_127; // @[ALU.scala 81:16 87:23]
  wire  _GEN_137 = 6'h2 == io_instr_id ? 1'h0 : _GEN_132; // @[ALU.scala 81:16 87:23]
  wire  _GEN_142 = 6'h1 == io_instr_id ? 1'h0 : _GEN_137; // @[ALU.scala 81:16 87:23]
  wire  branch_taken = 6'h0 == io_instr_id ? 1'h0 : _GEN_142; // @[ALU.scala 81:16 87:23]
  wire [31:0] _next_pc_T_11 = branch_taken ? _result_T_7 : _next_pc_T_1; // @[ALU.scala 126:21]
  wire [31:0] _GEN_0 = 6'h22 == io_instr_id | 6'h23 == io_instr_id | 6'h24 == io_instr_id ? _result_T_3 : 32'h0; // @[ALU.scala 156:14 80:10 87:23]
  wire [31:0] _GEN_2 = 6'h1d == io_instr_id | 6'h1e == io_instr_id | 6'h1f == io_instr_id | 6'h20 == io_instr_id | 6'h21
     == io_instr_id ? _result_T_3 : _GEN_0; // @[ALU.scala 151:14 87:23]
  wire  _GEN_4 = 6'h1d == io_instr_id | 6'h1e == io_instr_id | 6'h1f == io_instr_id | 6'h20 == io_instr_id | 6'h21 ==
    io_instr_id ? 1'h0 : 6'h22 == io_instr_id | 6'h23 == io_instr_id | 6'h24 == io_instr_id; // @[ALU.scala 84:12 87:23]
  wire [31:0] _GEN_6 = 6'h1c == io_instr_id ? _next_pc_T_11 : _next_pc_T_1; // @[ALU.scala 146:15 82:11 87:23]
  wire [31:0] _GEN_7 = 6'h1c == io_instr_id ? 32'h0 : _GEN_2; // @[ALU.scala 80:10 87:23]
  wire  _GEN_8 = 6'h1c == io_instr_id ? 1'h0 : 6'h1d == io_instr_id | 6'h1e == io_instr_id | 6'h1f == io_instr_id | 6'h20
     == io_instr_id | 6'h21 == io_instr_id; // @[ALU.scala 83:11 87:23]
  wire  _GEN_9 = 6'h1c == io_instr_id ? 1'h0 : _GEN_4; // @[ALU.scala 84:12 87:23]
  wire [31:0] _GEN_11 = 6'h1b == io_instr_id ? _next_pc_T_11 : _GEN_6; // @[ALU.scala 142:15 87:23]
  wire [31:0] _GEN_12 = 6'h1b == io_instr_id ? 32'h0 : _GEN_7; // @[ALU.scala 80:10 87:23]
  wire  _GEN_13 = 6'h1b == io_instr_id ? 1'h0 : _GEN_8; // @[ALU.scala 83:11 87:23]
  wire  _GEN_14 = 6'h1b == io_instr_id ? 1'h0 : _GEN_9; // @[ALU.scala 84:12 87:23]
  wire [31:0] _GEN_16 = 6'h1a == io_instr_id ? _next_pc_T_11 : _GEN_11; // @[ALU.scala 138:15 87:23]
  wire [31:0] _GEN_17 = 6'h1a == io_instr_id ? 32'h0 : _GEN_12; // @[ALU.scala 80:10 87:23]
  wire  _GEN_18 = 6'h1a == io_instr_id ? 1'h0 : _GEN_13; // @[ALU.scala 83:11 87:23]
  wire  _GEN_19 = 6'h1a == io_instr_id ? 1'h0 : _GEN_14; // @[ALU.scala 84:12 87:23]
  wire [31:0] _GEN_21 = 6'h19 == io_instr_id ? _next_pc_T_11 : _GEN_16; // @[ALU.scala 134:15 87:23]
  wire [31:0] _GEN_22 = 6'h19 == io_instr_id ? 32'h0 : _GEN_17; // @[ALU.scala 80:10 87:23]
  wire  _GEN_23 = 6'h19 == io_instr_id ? 1'h0 : _GEN_18; // @[ALU.scala 83:11 87:23]
  wire  _GEN_24 = 6'h19 == io_instr_id ? 1'h0 : _GEN_19; // @[ALU.scala 84:12 87:23]
  wire [31:0] _GEN_26 = 6'h18 == io_instr_id ? _next_pc_T_11 : _GEN_21; // @[ALU.scala 130:15 87:23]
  wire [31:0] _GEN_27 = 6'h18 == io_instr_id ? 32'h0 : _GEN_22; // @[ALU.scala 80:10 87:23]
  wire  _GEN_28 = 6'h18 == io_instr_id ? 1'h0 : _GEN_23; // @[ALU.scala 83:11 87:23]
  wire  _GEN_29 = 6'h18 == io_instr_id ? 1'h0 : _GEN_24; // @[ALU.scala 84:12 87:23]
  wire [31:0] _GEN_31 = 6'h17 == io_instr_id ? _next_pc_T_11 : _GEN_26; // @[ALU.scala 126:15 87:23]
  wire [31:0] _GEN_32 = 6'h17 == io_instr_id ? 32'h0 : _GEN_27; // @[ALU.scala 80:10 87:23]
  wire  _GEN_33 = 6'h17 == io_instr_id ? 1'h0 : _GEN_28; // @[ALU.scala 83:11 87:23]
  wire  _GEN_34 = 6'h17 == io_instr_id ? 1'h0 : _GEN_29; // @[ALU.scala 84:12 87:23]
  wire [31:0] _GEN_35 = 6'h16 == io_instr_id ? _next_pc_T_1 : _GEN_32; // @[ALU.scala 118:14 87:23]
  wire [31:0] _GEN_36 = 6'h16 == io_instr_id ? _next_pc_T_6 : _GEN_31; // @[ALU.scala 119:15 87:23]
  wire  _GEN_38 = 6'h16 == io_instr_id ? 1'h0 : _GEN_33; // @[ALU.scala 83:11 87:23]
  wire  _GEN_39 = 6'h16 == io_instr_id ? 1'h0 : _GEN_34; // @[ALU.scala 84:12 87:23]
  wire [31:0] _GEN_40 = 6'h15 == io_instr_id ? _next_pc_T_1 : _GEN_35; // @[ALU.scala 113:14 87:23]
  wire [31:0] _GEN_41 = 6'h15 == io_instr_id ? _result_T_7 : _GEN_36; // @[ALU.scala 114:15 87:23]
  wire  _GEN_43 = 6'h15 == io_instr_id ? 1'h0 : _GEN_38; // @[ALU.scala 83:11 87:23]
  wire  _GEN_44 = 6'h15 == io_instr_id ? 1'h0 : _GEN_39; // @[ALU.scala 84:12 87:23]
  wire [31:0] _GEN_45 = 6'h14 == io_instr_id ? {{31'd0}, io_src1_in < io_imm_in} : _GEN_40; // @[ALU.scala 87:23 109:24]
  wire [31:0] _GEN_46 = 6'h14 == io_instr_id ? _next_pc_T_1 : _GEN_41; // @[ALU.scala 82:11 87:23]
  wire  _GEN_48 = 6'h14 == io_instr_id ? 1'h0 : _GEN_43; // @[ALU.scala 83:11 87:23]
  wire  _GEN_49 = 6'h14 == io_instr_id ? 1'h0 : _GEN_44; // @[ALU.scala 84:12 87:23]
  wire [31:0] _GEN_50 = 6'h13 == io_instr_id ? {{31'd0}, io_src1_in < io_src2_in} : _GEN_45; // @[ALU.scala 87:23 108:24]
  wire [31:0] _GEN_51 = 6'h13 == io_instr_id ? _next_pc_T_1 : _GEN_46; // @[ALU.scala 82:11 87:23]
  wire  _GEN_53 = 6'h13 == io_instr_id ? 1'h0 : _GEN_48; // @[ALU.scala 83:11 87:23]
  wire  _GEN_54 = 6'h13 == io_instr_id ? 1'h0 : _GEN_49; // @[ALU.scala 84:12 87:23]
  wire [31:0] _GEN_55 = 6'h12 == io_instr_id ? {{31'd0}, $signed(_result_T_16) < $signed(_result_T_34)} : _GEN_50; // @[ALU.scala 87:23 107:24]
  wire [31:0] _GEN_56 = 6'h12 == io_instr_id ? _next_pc_T_1 : _GEN_51; // @[ALU.scala 82:11 87:23]
  wire  _GEN_58 = 6'h12 == io_instr_id ? 1'h0 : _GEN_53; // @[ALU.scala 83:11 87:23]
  wire  _GEN_59 = 6'h12 == io_instr_id ? 1'h0 : _GEN_54; // @[ALU.scala 84:12 87:23]
  wire [31:0] _GEN_60 = 6'h11 == io_instr_id ? {{31'd0}, $signed(_result_T_16) < $signed(_result_T_31)} : _GEN_55; // @[ALU.scala 87:23 106:24]
  wire [31:0] _GEN_61 = 6'h11 == io_instr_id ? _next_pc_T_1 : _GEN_56; // @[ALU.scala 82:11 87:23]
  wire  _GEN_63 = 6'h11 == io_instr_id ? 1'h0 : _GEN_58; // @[ALU.scala 83:11 87:23]
  wire  _GEN_64 = 6'h11 == io_instr_id ? 1'h0 : _GEN_59; // @[ALU.scala 84:12 87:23]
  wire [31:0] _GEN_65 = 6'h10 == io_instr_id ? _result_T_29 : _GEN_60; // @[ALU.scala 87:23 105:24]
  wire [31:0] _GEN_66 = 6'h10 == io_instr_id ? _next_pc_T_1 : _GEN_61; // @[ALU.scala 82:11 87:23]
  wire  _GEN_68 = 6'h10 == io_instr_id ? 1'h0 : _GEN_63; // @[ALU.scala 83:11 87:23]
  wire  _GEN_69 = 6'h10 == io_instr_id ? 1'h0 : _GEN_64; // @[ALU.scala 84:12 87:23]
  wire [31:0] _GEN_70 = 6'hf == io_instr_id ? _result_T_28 : _GEN_65; // @[ALU.scala 87:23 104:24]
  wire [31:0] _GEN_71 = 6'hf == io_instr_id ? _next_pc_T_1 : _GEN_66; // @[ALU.scala 82:11 87:23]
  wire  _GEN_73 = 6'hf == io_instr_id ? 1'h0 : _GEN_68; // @[ALU.scala 83:11 87:23]
  wire  _GEN_74 = 6'hf == io_instr_id ? 1'h0 : _GEN_69; // @[ALU.scala 84:12 87:23]
  wire [31:0] _GEN_75 = 6'he == io_instr_id ? _result_T_27 : _GEN_70; // @[ALU.scala 87:23 103:24]
  wire [31:0] _GEN_76 = 6'he == io_instr_id ? _next_pc_T_1 : _GEN_71; // @[ALU.scala 82:11 87:23]
  wire  _GEN_78 = 6'he == io_instr_id ? 1'h0 : _GEN_73; // @[ALU.scala 83:11 87:23]
  wire  _GEN_79 = 6'he == io_instr_id ? 1'h0 : _GEN_74; // @[ALU.scala 84:12 87:23]
  wire [31:0] _GEN_80 = 6'hd == io_instr_id ? _result_T_26 : _GEN_75; // @[ALU.scala 87:23 102:24]
  wire [31:0] _GEN_81 = 6'hd == io_instr_id ? _next_pc_T_1 : _GEN_76; // @[ALU.scala 82:11 87:23]
  wire  _GEN_83 = 6'hd == io_instr_id ? 1'h0 : _GEN_78; // @[ALU.scala 83:11 87:23]
  wire  _GEN_84 = 6'hd == io_instr_id ? 1'h0 : _GEN_79; // @[ALU.scala 84:12 87:23]
  wire [31:0] _GEN_85 = 6'hc == io_instr_id ? _result_T_25 : _GEN_80; // @[ALU.scala 87:23 101:24]
  wire [31:0] _GEN_86 = 6'hc == io_instr_id ? _next_pc_T_1 : _GEN_81; // @[ALU.scala 82:11 87:23]
  wire  _GEN_88 = 6'hc == io_instr_id ? 1'h0 : _GEN_83; // @[ALU.scala 83:11 87:23]
  wire  _GEN_89 = 6'hc == io_instr_id ? 1'h0 : _GEN_84; // @[ALU.scala 84:12 87:23]
  wire [31:0] _GEN_90 = 6'hb == io_instr_id ? _result_T_24 : _GEN_85; // @[ALU.scala 87:23 100:24]
  wire [31:0] _GEN_91 = 6'hb == io_instr_id ? _next_pc_T_1 : _GEN_86; // @[ALU.scala 82:11 87:23]
  wire  _GEN_93 = 6'hb == io_instr_id ? 1'h0 : _GEN_88; // @[ALU.scala 83:11 87:23]
  wire  _GEN_94 = 6'hb == io_instr_id ? 1'h0 : _GEN_89; // @[ALU.scala 84:12 87:23]
  wire [31:0] _GEN_95 = 6'ha == io_instr_id ? _result_T_23 : _GEN_90; // @[ALU.scala 87:23 99:24]
  wire [31:0] _GEN_96 = 6'ha == io_instr_id ? _next_pc_T_1 : _GEN_91; // @[ALU.scala 82:11 87:23]
  wire  _GEN_98 = 6'ha == io_instr_id ? 1'h0 : _GEN_93; // @[ALU.scala 83:11 87:23]
  wire  _GEN_99 = 6'ha == io_instr_id ? 1'h0 : _GEN_94; // @[ALU.scala 84:12 87:23]
  wire [31:0] _GEN_100 = 6'h9 == io_instr_id ? _result_T_19 : _GEN_95; // @[ALU.scala 87:23 98:24]
  wire [31:0] _GEN_101 = 6'h9 == io_instr_id ? _next_pc_T_1 : _GEN_96; // @[ALU.scala 82:11 87:23]
  wire  _GEN_103 = 6'h9 == io_instr_id ? 1'h0 : _GEN_98; // @[ALU.scala 83:11 87:23]
  wire  _GEN_104 = 6'h9 == io_instr_id ? 1'h0 : _GEN_99; // @[ALU.scala 84:12 87:23]
  wire [31:0] _GEN_105 = 6'h8 == io_instr_id ? _result_T_15 : _GEN_100; // @[ALU.scala 87:23 97:24]
  wire [31:0] _GEN_106 = 6'h8 == io_instr_id ? _next_pc_T_1 : _GEN_101; // @[ALU.scala 82:11 87:23]
  wire  _GEN_108 = 6'h8 == io_instr_id ? 1'h0 : _GEN_103; // @[ALU.scala 83:11 87:23]
  wire  _GEN_109 = 6'h8 == io_instr_id ? 1'h0 : _GEN_104; // @[ALU.scala 84:12 87:23]
  wire [31:0] _GEN_110 = 6'h7 == io_instr_id ? _result_T_13 : _GEN_105; // @[ALU.scala 87:23 96:24]
  wire [31:0] _GEN_111 = 6'h7 == io_instr_id ? _next_pc_T_1 : _GEN_106; // @[ALU.scala 82:11 87:23]
  wire  _GEN_113 = 6'h7 == io_instr_id ? 1'h0 : _GEN_108; // @[ALU.scala 83:11 87:23]
  wire  _GEN_114 = 6'h7 == io_instr_id ? 1'h0 : _GEN_109; // @[ALU.scala 84:12 87:23]
  wire [62:0] _GEN_115 = 6'h6 == io_instr_id ? _result_T_11 : {{31'd0}, _GEN_110}; // @[ALU.scala 87:23 95:24]
  wire [31:0] _GEN_116 = 6'h6 == io_instr_id ? _next_pc_T_1 : _GEN_111; // @[ALU.scala 82:11 87:23]
  wire  _GEN_118 = 6'h6 == io_instr_id ? 1'h0 : _GEN_113; // @[ALU.scala 83:11 87:23]
  wire  _GEN_119 = 6'h6 == io_instr_id ? 1'h0 : _GEN_114; // @[ALU.scala 84:12 87:23]
  wire [62:0] _GEN_120 = 6'h5 == io_instr_id ? _result_T_9 : _GEN_115; // @[ALU.scala 87:23 94:24]
  wire [31:0] _GEN_121 = 6'h5 == io_instr_id ? _next_pc_T_1 : _GEN_116; // @[ALU.scala 82:11 87:23]
  wire  _GEN_123 = 6'h5 == io_instr_id ? 1'h0 : _GEN_118; // @[ALU.scala 83:11 87:23]
  wire  _GEN_124 = 6'h5 == io_instr_id ? 1'h0 : _GEN_119; // @[ALU.scala 84:12 87:23]
  wire [62:0] _GEN_125 = 6'h4 == io_instr_id ? {{31'd0}, _result_T_7} : _GEN_120; // @[ALU.scala 87:23 93:24]
  wire [31:0] _GEN_126 = 6'h4 == io_instr_id ? _next_pc_T_1 : _GEN_121; // @[ALU.scala 82:11 87:23]
  wire  _GEN_128 = 6'h4 == io_instr_id ? 1'h0 : _GEN_123; // @[ALU.scala 83:11 87:23]
  wire  _GEN_129 = 6'h4 == io_instr_id ? 1'h0 : _GEN_124; // @[ALU.scala 84:12 87:23]
  wire [62:0] _GEN_130 = 6'h3 == io_instr_id ? {{31'd0}, io_imm_in} : _GEN_125; // @[ALU.scala 87:23 92:24]
  wire [31:0] _GEN_131 = 6'h3 == io_instr_id ? _next_pc_T_1 : _GEN_126; // @[ALU.scala 82:11 87:23]
  wire  _GEN_133 = 6'h3 == io_instr_id ? 1'h0 : _GEN_128; // @[ALU.scala 83:11 87:23]
  wire  _GEN_134 = 6'h3 == io_instr_id ? 1'h0 : _GEN_129; // @[ALU.scala 84:12 87:23]
  wire [62:0] _GEN_135 = 6'h2 == io_instr_id ? {{31'd0}, _result_T_5} : _GEN_130; // @[ALU.scala 87:23 91:24]
  wire [31:0] _GEN_136 = 6'h2 == io_instr_id ? _next_pc_T_1 : _GEN_131; // @[ALU.scala 82:11 87:23]
  wire  _GEN_138 = 6'h2 == io_instr_id ? 1'h0 : _GEN_133; // @[ALU.scala 83:11 87:23]
  wire  _GEN_139 = 6'h2 == io_instr_id ? 1'h0 : _GEN_134; // @[ALU.scala 84:12 87:23]
  wire [62:0] _GEN_140 = 6'h1 == io_instr_id ? {{31'd0}, _result_T_3} : _GEN_135; // @[ALU.scala 87:23 90:24]
  wire [31:0] _GEN_141 = 6'h1 == io_instr_id ? _next_pc_T_1 : _GEN_136; // @[ALU.scala 82:11 87:23]
  wire  _GEN_143 = 6'h1 == io_instr_id ? 1'h0 : _GEN_138; // @[ALU.scala 83:11 87:23]
  wire  _GEN_144 = 6'h1 == io_instr_id ? 1'h0 : _GEN_139; // @[ALU.scala 84:12 87:23]
  wire [62:0] _GEN_145 = 6'h0 == io_instr_id ? {{31'd0}, _result_T_1} : _GEN_140; // @[ALU.scala 87:23 89:24]
  wire [31:0] next_pc = 6'h0 == io_instr_id ? _next_pc_T_1 : _GEN_141; // @[ALU.scala 82:11 87:23]
  wire  is_load = 6'h0 == io_instr_id ? 1'h0 : _GEN_143; // @[ALU.scala 83:11 87:23]
  wire  is_store = 6'h0 == io_instr_id ? 1'h0 : _GEN_144; // @[ALU.scala 84:12 87:23]
  wire  valid = io_valid_in & ~io_flush_in; // @[ALU.scala 162:27]
  wire [31:0] result = _GEN_145[31:0]; // @[ALU.scala 73:20]
  wire  _io_branch_out_T = valid & branch_taken; // @[ALU.scala 165:26]
  assign io_result_out = valid ? result : 32'h0; // @[ALU.scala 163:23]
  assign io_valid_out = io_valid_in & ~io_flush_in; // @[ALU.scala 162:27]
  assign io_branch_out = valid & branch_taken; // @[ALU.scala 165:26]
  assign io_jump_addr = _io_branch_out_T ? next_pc : 32'h0; // @[ALU.scala 166:23]
  assign io_is_load = valid & is_load; // @[ALU.scala 167:26]
  assign io_is_store = valid & is_store; // @[ALU.scala 168:26]
endmodule
